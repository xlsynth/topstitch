// SPDX-License-Identifier: Apache-2.0

package pack;
    localparam int DefaultM = 8;
    localparam int DefaultN = 16;
endpackage
